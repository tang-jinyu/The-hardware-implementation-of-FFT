`timescale 1ns/1ps
module top#(
    parameter   N = 16,
    parameter   Q = 8
)
(
    input   clk2,
    input   rst,

    input   [N-1:0] in,
    output  [N-1:0] serial_out
);


    first_reg#(.N(N),.Q(Q))first_reg1
    (
        .clk2    (clk2),
        .rst     (rst ),
        .in      (in  ),
        .in0_r_0 (in0_r),
        .in1_r_0 (in1_r),
        .in2_r_0 (in2_r),
        .in3_r_0 (in3_r),
        .in4_r_0 (in4_r),
        .in5_r_0 (in5_r),
        .in6_r_0 (in6_r),
        .in7_r_0 (in7_r),
        .in8_r_0 (in8_r),
        .in9_r_0 (in9_r),
        .in10_r_0(in10_r),
        .in11_r_0(in11_r),
        .in12_r_0(in12_r),
        .in13_r_0(in13_r),
        .in14_r_0(in14_r),
        .in15_r_0(in15_r),
        .in16_r_0(in16_r),
        .in17_r_0(in17_r),
        .in18_r_0(in18_r),
        .in19_r_0(in19_r),
        .in20_r_0(in20_r),
        .in21_r_0(in21_r),
        .in22_r_0(in22_r),
        .in23_r_0(in23_r),
        .in24_r_0(in24_r),
        .in25_r_0(in25_r),
        .in26_r_0(in26_r),
        .in27_r_0(in27_r),
        .in28_r_0(in28_r),
        .in29_r_0(in29_r),
        .in30_r_0(in30_r),
        .in31_r_0(in31_r)
    );

    certain#(.N(N),.Q(Q)) certain1
    (
        .rst    (rst ),
        .clk2   (clk2),
        .in0_r  (in0_r),
        .in1_r  (in1_r),
        .in2_r  (in2_r),
        .in3_r  (in3_r),
        .in4_r  (in4_r),
        .in5_r  (in5_r),
        .in6_r  (in6_r),
        .in7_r  (in7_r),
        .in8_r  (in8_r),
        .in9_r  (in9_r),
        .in10_r (in10_r),
        .in11_r (in11_r),
        .in12_r (in12_r),
        .in13_r (in13_r),
        .in14_r (in14_r),
        .in15_r (in15_r),
        .in16_r (in16_r),
        .in17_r (in17_r),
        .in18_r (in18_r),
        .in19_r (in19_r),
        .in20_r (in20_r),
        .in21_r (in21_r),
        .in22_r (in22_r),
        .in23_r (in23_r),
        .in24_r (in24_r),
        .in25_r (in25_r),
        .in26_r (in26_r),
        .in27_r (in27_r),
        .in28_r (in28_r),
        .in29_r (in29_r),
        .in30_r (in30_r),
        .in31_r (in31_r),

        .out0_r (out0_r ),
        .out1_r (out1_r ),
        .out2_r (out2_r ),
        .out3_r (out3_r ),
        .out4_r (out4_r ),
        .out5_r (out5_r ),
        .out6_r (out6_r ),
        .out7_r (out7_r ),
        .out8_r (out8_r ),
        .out9_r (out9_r ),
        .out10_r(out10_r),
        .out11_r(out11_r),
        .out12_r(out12_r),
        .out13_r(out13_r),
        .out14_r(out14_r),
        .out15_r(out15_r),
        .out16_r(out16_r),
        .out17_r(out17_r),
        .out18_r(out18_r),
        .out19_r(out19_r),
        .out20_r(out20_r),
        .out21_r(out21_r),
        .out22_r(out22_r),
        .out23_r(out23_r),
        .out24_r(out24_r),
        .out25_r(out25_r),
        .out26_r(out26_r),
        .out27_r(out27_r),
        .out28_r(out28_r),
        .out29_r(out29_r),
        .out30_r(out30_r),
        .out31_r(out31_r),
        
        .out0_i (out0_i ),
        .out1_i (out1_i ),
        .out2_i (out2_i ),
        .out3_i (out3_i ),
        .out4_i (out4_i ),
        .out5_i (out5_i ),
        .out6_i (out6_i ),
        .out7_i (out7_i ),
        .out8_i (out8_i ),
        .out9_i (out9_i ),
        .out10_i(out10_i),
        .out11_i(out11_i),
        .out12_i(out12_i),
        .out13_i(out13_i),
        .out14_i(out14_i),
        .out15_i(out15_i),
        .out16_i(out16_i),
        .out17_i(out17_i),
        .out18_i(out18_i),
        .out19_i(out19_i),
        .out20_i(out20_i),
        .out21_i(out21_i),
        .out22_i(out22_i),
        .out23_i(out23_i),
        .out24_i(out24_i),
        .out25_i(out25_i),
        .out26_i(out26_i),
        .out27_i(out27_i),
        .out28_i(out28_i),
        .out29_i(out29_i),
        .out30_i(out30_i),
        .out31_i(out31_i)
    );

    post_reg#(.N(N),.Q(Q))post_reg1
    (
        .clk2           (clk2),
        .rst            (rst ),
        .out0_r         (out0_r),
        .out0_i         (out0_i),
        .out1_r         (out1_r),
        .out1_i         (out1_i),
        .out2_r         (out2_r),
        .out2_i         (out2_i),
        .out3_r         (out3_r),
        .out3_i         (out3_i),
        .out4_r         (out4_r),
        .out4_i         (out4_i),
        .out5_r         (out5_r),
        .out5_i         (out5_i),
        .out6_r         (out6_r),
        .out6_i         (out6_i),
        .out7_r         (out7_r),
        .out7_i         (out7_i),
        .out8_r         (out8_r),
        .out8_i         (out8_i),
        .out9_r         (out9_r),
        .out9_i         (out9_i),
        .out10_r        (out10_r),
        .out10_i        (out10_i),
        .out11_r        (out11_r),
        .out11_i        (out11_i),
        .out12_r        (out12_r),
        .out12_i        (out12_i),
        .out13_r        (out13_r),
        .out13_i        (out13_i),
        .out14_r        (out14_r),
        .out14_i        (out14_i),
        .out15_r        (out15_r),
        .out15_i        (out15_i),
        .out16_r        (out16_r),
        .out16_i        (out16_i),
        .out17_r        (out17_r),
        .out17_i        (out17_i),
        .out18_r        (out18_r),
        .out18_i        (out18_i),
        .out19_r        (out19_r),
        .out19_i        (out19_i),
        .out20_r        (out20_r),
        .out20_i        (out20_i),
        .out21_r        (out21_r),
        .out21_i        (out21_i),
        .out22_r        (out22_r),
        .out22_i        (out22_i),
        .out23_r        (out23_r),
        .out23_i        (out23_i),
        .out24_r        (out24_r),
        .out24_i        (out24_i),
        .out25_r        (out25_r),
        .out25_i        (out25_i),
        .out26_r        (out26_r),
        .out26_i        (out26_i),
        .out27_r        (out27_r),
        .out27_i        (out27_i),
        .out28_r        (out28_r),
        .out28_i        (out28_i),
        .out29_r        (out29_r),
        .out29_i        (out29_i),
        .out30_r        (out30_r),
        .out30_i        (out30_i),
        .out31_r        (out31_r),
        .out31_i        (out31_i),
        .serial_out     (serial_out ),
        .out_valid      (out_valid),
        .out_type       (out_type   ),
        .output_busy    (output_busy),
        .output_done    (output_done)
    );
endmodule